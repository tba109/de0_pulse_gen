//////////////////////////////////////////////////////////////////////////////////////
// Tyler Anderson Wed Dec  5 16:41:30 EST 2018
// exp_pgen.v
//
//////////////////////////////////////////////////////////////////////////////////////
module exp_pgen
  (
   
   );

endmodule
