module version_number
  (
   output [15:0] vnum
   );

   assign vnum = 16'd1;

endmodule
  
