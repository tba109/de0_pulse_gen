///////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Tyler Anderson Tue Aug 14 17:13:35 EDT 2018
//
// gaus_rand_tb.v
//
// Gaussian Random number generator
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////

`timescale 1ns/1ns

///////////////////////////////////////////////////////////////////////////////////////////////////
// Test cases
///////////////////////////////////////////////////////////////////////////////////////////////////
`define TEST_CASE_SIMPLE

module gaus_rand_tb;
   
   //////////////////////////////////////////////////////////////////////
   // I/O
   //////////////////////////////////////////////////////////////////////   
   parameter SYSCLK_PERIOD = 10;
   reg clk;
   reg rst;
   wire [11:0] gr;
   integer     fout; 
   
   // Connections
   
   //////////////////////////////////////////////////////////////////////
   // Clock Driver
   //////////////////////////////////////////////////////////////////////
   always @(clk)
     #(SYSCLK_PERIOD / 2.0) clk <= !clk;
				   
   //////////////////////////////////////////////////////////////////////
   // Simulated interfaces
   //////////////////////////////////////////////////////////////////////   
      
   //////////////////////////////////////////////////////////////////////
   // UUT
   //////////////////////////////////////////////////////////////////////   
   gaus_rand GR_0(.clk(clk),.gr(gr)); 
   
   //////////////////////////////////////////////////////////////////////
   // Test case
   //////////////////////////////////////////////////////////////////////   
   `ifdef TEST_CASE_SIMPLE
   
   initial
     begin
	// fout = $fopen("gr.txt","w"); 
	clk <= 0;
	rst <= 1; 
	// Reset	
	#(10 * SYSCLK_PERIOD);
	rst <= 1'b0;

	// Logging
	$display("");
	$display("------------------------------------------------------");
	$display("Test Case: TEST_CASE_SIMPLE");

	#(100_000); 
	
	// $fclose(fout);
	// Stimulate UUT
     end
   // always @(posedge clk) $write(fout,"%x\n",gr);
   always @(posedge clk) $display("%03x",gr); 
   `endif

   //////////////////////////////////////////////////////////////////////
   // Tasks (e.g., writing data, etc.)
   //////////////////////////////////////////////////////////////////////   
   
   
   
endmodule

// Local Variables:
// verilog-library-flags:("-y ../hdl/")
// End:
   
