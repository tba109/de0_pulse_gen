// DE0_CV_system.v

// Generated using ACDS version 14.0 209 at 2014.11.17.10:01:09

`timescale 1 ps / 1 ps
module DE0_CV_system (
		input  wire       clk_clk,                                //                             clk.clk
		output wire       sd_clk_export,                          //                          sd_clk.export
		inout  wire       sd_cmd_export,                          //                          sd_cmd.export
		inout  wire [3:0] sd_dat_export,                          //                          sd_dat.export
		output wire [9:0] ledr_external_connection_export,        //        ledr_external_connection.export
		input  wire [3:0] key_external_connection_export,         //         key_external_connection.export
		input  wire       cpu_reset_n_external_connection_export, // cpu_reset_n_external_connection.export
		input  wire       reset_reset_n                           //                           reset.reset_n
	);

	wire         pll_100_outclk0_clk;                                         // pll_100:outclk_0 -> [cpu:clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, irq_synchronizer_002:sender_clk, irq_synchronizer_003:sender_clk, mm_clock_crossing_bridge:s0_clk, mm_interconnect_0:pll_100_outclk0_clk, onchip_memory:clk, rst_controller:clk, rst_controller_002:clk]
	wire         cpu_instruction_master_waitrequest;                          // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [19:0] cpu_instruction_master_address;                              // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                 // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire  [31:0] cpu_instruction_master_readdata;                             // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_readdatavalid;                        // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire         cpu_data_master_waitrequest;                                 // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire  [31:0] cpu_data_master_writedata;                                   // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [24:0] cpu_data_master_address;                                     // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire         cpu_data_master_write;                                       // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire         cpu_data_master_read;                                        // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire  [31:0] cpu_data_master_readdata;                                    // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_debugaccess;                                 // cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire         cpu_data_master_readdatavalid;                               // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire   [3:0] cpu_data_master_byteenable;                                  // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;         // cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;           // mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;             // mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;               // mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;                // mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;            // cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;         // mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;          // mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;                // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire  [14:0] mm_interconnect_0_onchip_memory_s1_address;                  // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;               // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire         mm_interconnect_0_onchip_memory_s1_clken;                    // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire         mm_interconnect_0_onchip_memory_s1_write;                    // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;                 // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;               // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;   // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;    // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;      // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_waitrequest;   // mm_clock_crossing_bridge:s0_waitrequest -> mm_interconnect_0:mm_clock_crossing_bridge_s0_waitrequest
	wire   [0:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_burstcount;    // mm_interconnect_0:mm_clock_crossing_bridge_s0_burstcount -> mm_clock_crossing_bridge:s0_burstcount
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_writedata;     // mm_interconnect_0:mm_clock_crossing_bridge_s0_writedata -> mm_clock_crossing_bridge:s0_writedata
	wire  [11:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_address;       // mm_interconnect_0:mm_clock_crossing_bridge_s0_address -> mm_clock_crossing_bridge:s0_address
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_write;         // mm_interconnect_0:mm_clock_crossing_bridge_s0_write -> mm_clock_crossing_bridge:s0_write
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_read;          // mm_interconnect_0:mm_clock_crossing_bridge_s0_read -> mm_clock_crossing_bridge:s0_read
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_readdata;      // mm_clock_crossing_bridge:s0_readdata -> mm_interconnect_0:mm_clock_crossing_bridge_s0_readdata
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_debugaccess;   // mm_interconnect_0:mm_clock_crossing_bridge_s0_debugaccess -> mm_clock_crossing_bridge:s0_debugaccess
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_readdatavalid; // mm_clock_crossing_bridge:s0_readdatavalid -> mm_interconnect_0:mm_clock_crossing_bridge_s0_readdatavalid
	wire   [3:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_byteenable;    // mm_interconnect_0:mm_clock_crossing_bridge_s0_byteenable -> mm_clock_crossing_bridge:s0_byteenable
	wire   [0:0] mm_clock_crossing_bridge_m0_burstcount;                      // mm_clock_crossing_bridge:m0_burstcount -> mm_interconnect_1:mm_clock_crossing_bridge_m0_burstcount
	wire         mm_clock_crossing_bridge_m0_waitrequest;                     // mm_interconnect_1:mm_clock_crossing_bridge_m0_waitrequest -> mm_clock_crossing_bridge:m0_waitrequest
	wire  [11:0] mm_clock_crossing_bridge_m0_address;                         // mm_clock_crossing_bridge:m0_address -> mm_interconnect_1:mm_clock_crossing_bridge_m0_address
	wire  [31:0] mm_clock_crossing_bridge_m0_writedata;                       // mm_clock_crossing_bridge:m0_writedata -> mm_interconnect_1:mm_clock_crossing_bridge_m0_writedata
	wire         mm_clock_crossing_bridge_m0_write;                           // mm_clock_crossing_bridge:m0_write -> mm_interconnect_1:mm_clock_crossing_bridge_m0_write
	wire         mm_clock_crossing_bridge_m0_read;                            // mm_clock_crossing_bridge:m0_read -> mm_interconnect_1:mm_clock_crossing_bridge_m0_read
	wire  [31:0] mm_clock_crossing_bridge_m0_readdata;                        // mm_interconnect_1:mm_clock_crossing_bridge_m0_readdata -> mm_clock_crossing_bridge:m0_readdata
	wire         mm_clock_crossing_bridge_m0_debugaccess;                     // mm_clock_crossing_bridge:m0_debugaccess -> mm_interconnect_1:mm_clock_crossing_bridge_m0_debugaccess
	wire   [3:0] mm_clock_crossing_bridge_m0_byteenable;                      // mm_clock_crossing_bridge:m0_byteenable -> mm_interconnect_1:mm_clock_crossing_bridge_m0_byteenable
	wire         mm_clock_crossing_bridge_m0_readdatavalid;                   // mm_interconnect_1:mm_clock_crossing_bridge_m0_readdatavalid -> mm_clock_crossing_bridge:m0_readdatavalid
	wire  [31:0] mm_interconnect_1_sd_clk_s1_writedata;                       // mm_interconnect_1:sd_clk_s1_writedata -> sd_clk:writedata
	wire   [1:0] mm_interconnect_1_sd_clk_s1_address;                         // mm_interconnect_1:sd_clk_s1_address -> sd_clk:address
	wire         mm_interconnect_1_sd_clk_s1_chipselect;                      // mm_interconnect_1:sd_clk_s1_chipselect -> sd_clk:chipselect
	wire         mm_interconnect_1_sd_clk_s1_write;                           // mm_interconnect_1:sd_clk_s1_write -> sd_clk:write_n
	wire  [31:0] mm_interconnect_1_sd_clk_s1_readdata;                        // sd_clk:readdata -> mm_interconnect_1:sd_clk_s1_readdata
	wire  [31:0] mm_interconnect_1_sd_cmd_s1_writedata;                       // mm_interconnect_1:sd_cmd_s1_writedata -> sd_cmd:writedata
	wire   [1:0] mm_interconnect_1_sd_cmd_s1_address;                         // mm_interconnect_1:sd_cmd_s1_address -> sd_cmd:address
	wire         mm_interconnect_1_sd_cmd_s1_chipselect;                      // mm_interconnect_1:sd_cmd_s1_chipselect -> sd_cmd:chipselect
	wire         mm_interconnect_1_sd_cmd_s1_write;                           // mm_interconnect_1:sd_cmd_s1_write -> sd_cmd:write_n
	wire  [31:0] mm_interconnect_1_sd_cmd_s1_readdata;                        // sd_cmd:readdata -> mm_interconnect_1:sd_cmd_s1_readdata
	wire  [31:0] mm_interconnect_1_sd_dat_s1_writedata;                       // mm_interconnect_1:sd_dat_s1_writedata -> sd_dat:writedata
	wire   [1:0] mm_interconnect_1_sd_dat_s1_address;                         // mm_interconnect_1:sd_dat_s1_address -> sd_dat:address
	wire         mm_interconnect_1_sd_dat_s1_chipselect;                      // mm_interconnect_1:sd_dat_s1_chipselect -> sd_dat:chipselect
	wire         mm_interconnect_1_sd_dat_s1_write;                           // mm_interconnect_1:sd_dat_s1_write -> sd_dat:write_n
	wire  [31:0] mm_interconnect_1_sd_dat_s1_readdata;                        // sd_dat:readdata -> mm_interconnect_1:sd_dat_s1_readdata
	wire  [31:0] mm_interconnect_1_ledr_s1_writedata;                         // mm_interconnect_1:ledr_s1_writedata -> ledr:writedata
	wire   [1:0] mm_interconnect_1_ledr_s1_address;                           // mm_interconnect_1:ledr_s1_address -> ledr:address
	wire         mm_interconnect_1_ledr_s1_chipselect;                        // mm_interconnect_1:ledr_s1_chipselect -> ledr:chipselect
	wire         mm_interconnect_1_ledr_s1_write;                             // mm_interconnect_1:ledr_s1_write -> ledr:write_n
	wire  [31:0] mm_interconnect_1_ledr_s1_readdata;                          // ledr:readdata -> mm_interconnect_1:ledr_s1_readdata
	wire  [31:0] mm_interconnect_1_key_s1_writedata;                          // mm_interconnect_1:key_s1_writedata -> key:writedata
	wire   [1:0] mm_interconnect_1_key_s1_address;                            // mm_interconnect_1:key_s1_address -> key:address
	wire         mm_interconnect_1_key_s1_chipselect;                         // mm_interconnect_1:key_s1_chipselect -> key:chipselect
	wire         mm_interconnect_1_key_s1_write;                              // mm_interconnect_1:key_s1_write -> key:write_n
	wire  [31:0] mm_interconnect_1_key_s1_readdata;                           // key:readdata -> mm_interconnect_1:key_s1_readdata
	wire  [31:0] mm_interconnect_1_cpu_reset_n_s1_writedata;                  // mm_interconnect_1:cpu_reset_n_s1_writedata -> cpu_reset_n:writedata
	wire   [1:0] mm_interconnect_1_cpu_reset_n_s1_address;                    // mm_interconnect_1:cpu_reset_n_s1_address -> cpu_reset_n:address
	wire         mm_interconnect_1_cpu_reset_n_s1_chipselect;                 // mm_interconnect_1:cpu_reset_n_s1_chipselect -> cpu_reset_n:chipselect
	wire         mm_interconnect_1_cpu_reset_n_s1_write;                      // mm_interconnect_1:cpu_reset_n_s1_write -> cpu_reset_n:write_n
	wire  [31:0] mm_interconnect_1_cpu_reset_n_s1_readdata;                   // cpu_reset_n:readdata -> mm_interconnect_1:cpu_reset_n_s1_readdata
	wire  [15:0] mm_interconnect_1_timer_1_s1_writedata;                      // mm_interconnect_1:timer_1_s1_writedata -> timer_1:writedata
	wire   [2:0] mm_interconnect_1_timer_1_s1_address;                        // mm_interconnect_1:timer_1_s1_address -> timer_1:address
	wire         mm_interconnect_1_timer_1_s1_chipselect;                     // mm_interconnect_1:timer_1_s1_chipselect -> timer_1:chipselect
	wire         mm_interconnect_1_timer_1_s1_write;                          // mm_interconnect_1:timer_1_s1_write -> timer_1:write_n
	wire  [15:0] mm_interconnect_1_timer_1_s1_readdata;                       // timer_1:readdata -> mm_interconnect_1:timer_1_s1_readdata
	wire  [31:0] cpu_d_irq_irq;                                               // irq_mapper:sender_irq -> cpu:d_irq
	wire         irq_mapper_receiver0_irq;                                    // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                               // key:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver1_irq;                                    // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                           // cpu_reset_n:irq -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_receiver2_irq;                                    // irq_synchronizer_002:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                           // timer_1:irq -> irq_synchronizer_002:receiver_irq
	wire         irq_mapper_receiver3_irq;                                    // irq_synchronizer_003:sender_irq -> irq_mapper:receiver3_irq
	wire   [0:0] irq_synchronizer_003_receiver_irq;                           // jtag_uart:av_irq -> irq_synchronizer_003:receiver_irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [cpu:reset_n, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, onchip_memory:reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [cpu:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	wire         cpu_jtag_debug_module_reset_reset;                           // cpu:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_003:reset_in1]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [cpu_reset_n:reset_n, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, key:reset_n, ledr:reset_n, mm_clock_crossing_bridge:m0_reset, mm_interconnect_1:mm_clock_crossing_bridge_m0_reset_reset_bridge_in_reset_reset, pll_100:rst, sd_clk:reset_n, sd_cmd:reset_n, sd_dat:reset_n, timer_1:reset_n]
	wire         rst_controller_002_reset_out_reset;                          // rst_controller_002:reset_out -> [mm_clock_crossing_bridge:s0_reset, mm_interconnect_0:mm_clock_crossing_bridge_s0_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_003_reset_out_reset;                          // rst_controller_003:reset_out -> [irq_synchronizer_003:receiver_reset, jtag_uart:rst_n, mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset]

	DE0_CV_system_cpu cpu (
		.clk                                   (pll_100_outclk0_clk),                                 //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                     //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (cpu_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	DE0_CV_system_sd_dat sd_dat (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_1_sd_dat_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_sd_dat_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_sd_dat_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_sd_dat_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_sd_dat_s1_readdata),   //                    .readdata
		.bidir_port (sd_dat_export)                           // external_connection.export
	);

	DE0_CV_system_sd_cmd sd_cmd (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_1_sd_cmd_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_sd_cmd_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_sd_cmd_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_sd_cmd_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_sd_cmd_s1_readdata),   //                    .readdata
		.bidir_port (sd_cmd_export)                           // external_connection.export
	);

	DE0_CV_system_sd_clk sd_clk (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_1_sd_clk_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_sd_clk_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_sd_clk_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_sd_clk_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_sd_clk_s1_readdata),   //                    .readdata
		.out_port   (sd_clk_export)                           // external_connection.export
	);

	DE0_CV_system_onchip_memory onchip_memory (
		.clk        (pll_100_outclk0_clk),                           //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)             //       .reset_req
	);

	DE0_CV_system_pll_100 pll_100 (
		.refclk   (clk_clk),                            //  refclk.clk
		.rst      (rst_controller_001_reset_out_reset), //   reset.reset
		.outclk_0 (pll_100_outclk0_clk),                // outclk0.clk
		.locked   ()                                    // (terminated)
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (12),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (4),
		.RESPONSE_FIFO_DEPTH (4),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) mm_clock_crossing_bridge (
		.m0_clk           (clk_clk),                                                     //   m0_clk.clk
		.m0_reset         (rst_controller_001_reset_out_reset),                          // m0_reset.reset
		.s0_clk           (pll_100_outclk0_clk),                                         //   s0_clk.clk
		.s0_reset         (rst_controller_002_reset_out_reset),                          // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_clock_crossing_bridge_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_clock_crossing_bridge_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_clock_crossing_bridge_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_clock_crossing_bridge_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_mm_clock_crossing_bridge_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_mm_clock_crossing_bridge_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_mm_clock_crossing_bridge_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_mm_clock_crossing_bridge_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_mm_clock_crossing_bridge_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_clock_crossing_bridge_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (mm_clock_crossing_bridge_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (mm_clock_crossing_bridge_m0_readdata),                        //         .readdata
		.m0_readdatavalid (mm_clock_crossing_bridge_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (mm_clock_crossing_bridge_m0_burstcount),                      //         .burstcount
		.m0_writedata     (mm_clock_crossing_bridge_m0_writedata),                       //         .writedata
		.m0_address       (mm_clock_crossing_bridge_m0_address),                         //         .address
		.m0_write         (mm_clock_crossing_bridge_m0_write),                           //         .write
		.m0_read          (mm_clock_crossing_bridge_m0_read),                            //         .read
		.m0_byteenable    (mm_clock_crossing_bridge_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (mm_clock_crossing_bridge_m0_debugaccess)                      //         .debugaccess
	);

	DE0_CV_system_ledr ledr (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_1_ledr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_ledr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_ledr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_ledr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_ledr_s1_readdata),   //                    .readdata
		.out_port   (ledr_external_connection_export)       // external_connection.export
	);

	DE0_CV_system_key key (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_1_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_key_s1_readdata),   //                    .readdata
		.in_port    (key_external_connection_export),      // external_connection.export
		.irq        (irq_synchronizer_receiver_irq)        //                 irq.irq
	);

	DE0_CV_system_cpu_reset_n cpu_reset_n (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_1_cpu_reset_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_cpu_reset_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_cpu_reset_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_cpu_reset_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_cpu_reset_n_s1_readdata),   //                    .readdata
		.in_port    (cpu_reset_n_external_connection_export),      // external_connection.export
		.irq        (irq_synchronizer_001_receiver_irq)            //                 irq.irq
	);

	DE0_CV_system_timer_1 timer_1 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_1_timer_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_1_s1_write),     //      .write_n
		.irq        (irq_synchronizer_002_receiver_irq)        //   irq.irq
	);

	DE0_CV_system_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_003_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_synchronizer_003_receiver_irq)                          //               irq.irq
	);

	DE0_CV_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                                 (clk_clk),                                                     //                                               clk_0_clk.clk
		.pll_100_outclk0_clk                                           (pll_100_outclk0_clk),                                         //                                         pll_100_outclk0.clk
		.cpu_reset_n_reset_bridge_in_reset_reset                       (rst_controller_reset_out_reset),                              //                       cpu_reset_n_reset_bridge_in_reset.reset
		.jtag_uart_reset_reset_bridge_in_reset_reset                   (rst_controller_003_reset_out_reset),                          //                   jtag_uart_reset_reset_bridge_in_reset.reset
		.mm_clock_crossing_bridge_s0_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                          // mm_clock_crossing_bridge_s0_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                                       (cpu_data_master_address),                                     //                                         cpu_data_master.address
		.cpu_data_master_waitrequest                                   (cpu_data_master_waitrequest),                                 //                                                        .waitrequest
		.cpu_data_master_byteenable                                    (cpu_data_master_byteenable),                                  //                                                        .byteenable
		.cpu_data_master_read                                          (cpu_data_master_read),                                        //                                                        .read
		.cpu_data_master_readdata                                      (cpu_data_master_readdata),                                    //                                                        .readdata
		.cpu_data_master_readdatavalid                                 (cpu_data_master_readdatavalid),                               //                                                        .readdatavalid
		.cpu_data_master_write                                         (cpu_data_master_write),                                       //                                                        .write
		.cpu_data_master_writedata                                     (cpu_data_master_writedata),                                   //                                                        .writedata
		.cpu_data_master_debugaccess                                   (cpu_data_master_debugaccess),                                 //                                                        .debugaccess
		.cpu_instruction_master_address                                (cpu_instruction_master_address),                              //                                  cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                            (cpu_instruction_master_waitrequest),                          //                                                        .waitrequest
		.cpu_instruction_master_read                                   (cpu_instruction_master_read),                                 //                                                        .read
		.cpu_instruction_master_readdata                               (cpu_instruction_master_readdata),                             //                                                        .readdata
		.cpu_instruction_master_readdatavalid                          (cpu_instruction_master_readdatavalid),                        //                                                        .readdatavalid
		.cpu_jtag_debug_module_address                                 (mm_interconnect_0_cpu_jtag_debug_module_address),             //                                   cpu_jtag_debug_module.address
		.cpu_jtag_debug_module_write                                   (mm_interconnect_0_cpu_jtag_debug_module_write),               //                                                        .write
		.cpu_jtag_debug_module_read                                    (mm_interconnect_0_cpu_jtag_debug_module_read),                //                                                        .read
		.cpu_jtag_debug_module_readdata                                (mm_interconnect_0_cpu_jtag_debug_module_readdata),            //                                                        .readdata
		.cpu_jtag_debug_module_writedata                               (mm_interconnect_0_cpu_jtag_debug_module_writedata),           //                                                        .writedata
		.cpu_jtag_debug_module_byteenable                              (mm_interconnect_0_cpu_jtag_debug_module_byteenable),          //                                                        .byteenable
		.cpu_jtag_debug_module_waitrequest                             (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),         //                                                        .waitrequest
		.cpu_jtag_debug_module_debugaccess                             (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),         //                                                        .debugaccess
		.jtag_uart_avalon_jtag_slave_address                           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),       //                             jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),         //                                                        .write
		.jtag_uart_avalon_jtag_slave_read                              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),          //                                                        .read
		.jtag_uart_avalon_jtag_slave_readdata                          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),      //                                                        .readdata
		.jtag_uart_avalon_jtag_slave_writedata                         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),     //                                                        .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),   //                                                        .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),    //                                                        .chipselect
		.mm_clock_crossing_bridge_s0_address                           (mm_interconnect_0_mm_clock_crossing_bridge_s0_address),       //                             mm_clock_crossing_bridge_s0.address
		.mm_clock_crossing_bridge_s0_write                             (mm_interconnect_0_mm_clock_crossing_bridge_s0_write),         //                                                        .write
		.mm_clock_crossing_bridge_s0_read                              (mm_interconnect_0_mm_clock_crossing_bridge_s0_read),          //                                                        .read
		.mm_clock_crossing_bridge_s0_readdata                          (mm_interconnect_0_mm_clock_crossing_bridge_s0_readdata),      //                                                        .readdata
		.mm_clock_crossing_bridge_s0_writedata                         (mm_interconnect_0_mm_clock_crossing_bridge_s0_writedata),     //                                                        .writedata
		.mm_clock_crossing_bridge_s0_burstcount                        (mm_interconnect_0_mm_clock_crossing_bridge_s0_burstcount),    //                                                        .burstcount
		.mm_clock_crossing_bridge_s0_byteenable                        (mm_interconnect_0_mm_clock_crossing_bridge_s0_byteenable),    //                                                        .byteenable
		.mm_clock_crossing_bridge_s0_readdatavalid                     (mm_interconnect_0_mm_clock_crossing_bridge_s0_readdatavalid), //                                                        .readdatavalid
		.mm_clock_crossing_bridge_s0_waitrequest                       (mm_interconnect_0_mm_clock_crossing_bridge_s0_waitrequest),   //                                                        .waitrequest
		.mm_clock_crossing_bridge_s0_debugaccess                       (mm_interconnect_0_mm_clock_crossing_bridge_s0_debugaccess),   //                                                        .debugaccess
		.onchip_memory_s1_address                                      (mm_interconnect_0_onchip_memory_s1_address),                  //                                        onchip_memory_s1.address
		.onchip_memory_s1_write                                        (mm_interconnect_0_onchip_memory_s1_write),                    //                                                        .write
		.onchip_memory_s1_readdata                                     (mm_interconnect_0_onchip_memory_s1_readdata),                 //                                                        .readdata
		.onchip_memory_s1_writedata                                    (mm_interconnect_0_onchip_memory_s1_writedata),                //                                                        .writedata
		.onchip_memory_s1_byteenable                                   (mm_interconnect_0_onchip_memory_s1_byteenable),               //                                                        .byteenable
		.onchip_memory_s1_chipselect                                   (mm_interconnect_0_onchip_memory_s1_chipselect),               //                                                        .chipselect
		.onchip_memory_s1_clken                                        (mm_interconnect_0_onchip_memory_s1_clken)                     //                                                        .clken
	);

	DE0_CV_system_mm_interconnect_1 mm_interconnect_1 (
		.clk_0_clk_clk                                                 (clk_clk),                                     //                                               clk_0_clk.clk
		.mm_clock_crossing_bridge_m0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),          // mm_clock_crossing_bridge_m0_reset_reset_bridge_in_reset.reset
		.mm_clock_crossing_bridge_m0_address                           (mm_clock_crossing_bridge_m0_address),         //                             mm_clock_crossing_bridge_m0.address
		.mm_clock_crossing_bridge_m0_waitrequest                       (mm_clock_crossing_bridge_m0_waitrequest),     //                                                        .waitrequest
		.mm_clock_crossing_bridge_m0_burstcount                        (mm_clock_crossing_bridge_m0_burstcount),      //                                                        .burstcount
		.mm_clock_crossing_bridge_m0_byteenable                        (mm_clock_crossing_bridge_m0_byteenable),      //                                                        .byteenable
		.mm_clock_crossing_bridge_m0_read                              (mm_clock_crossing_bridge_m0_read),            //                                                        .read
		.mm_clock_crossing_bridge_m0_readdata                          (mm_clock_crossing_bridge_m0_readdata),        //                                                        .readdata
		.mm_clock_crossing_bridge_m0_readdatavalid                     (mm_clock_crossing_bridge_m0_readdatavalid),   //                                                        .readdatavalid
		.mm_clock_crossing_bridge_m0_write                             (mm_clock_crossing_bridge_m0_write),           //                                                        .write
		.mm_clock_crossing_bridge_m0_writedata                         (mm_clock_crossing_bridge_m0_writedata),       //                                                        .writedata
		.mm_clock_crossing_bridge_m0_debugaccess                       (mm_clock_crossing_bridge_m0_debugaccess),     //                                                        .debugaccess
		.cpu_reset_n_s1_address                                        (mm_interconnect_1_cpu_reset_n_s1_address),    //                                          cpu_reset_n_s1.address
		.cpu_reset_n_s1_write                                          (mm_interconnect_1_cpu_reset_n_s1_write),      //                                                        .write
		.cpu_reset_n_s1_readdata                                       (mm_interconnect_1_cpu_reset_n_s1_readdata),   //                                                        .readdata
		.cpu_reset_n_s1_writedata                                      (mm_interconnect_1_cpu_reset_n_s1_writedata),  //                                                        .writedata
		.cpu_reset_n_s1_chipselect                                     (mm_interconnect_1_cpu_reset_n_s1_chipselect), //                                                        .chipselect
		.key_s1_address                                                (mm_interconnect_1_key_s1_address),            //                                                  key_s1.address
		.key_s1_write                                                  (mm_interconnect_1_key_s1_write),              //                                                        .write
		.key_s1_readdata                                               (mm_interconnect_1_key_s1_readdata),           //                                                        .readdata
		.key_s1_writedata                                              (mm_interconnect_1_key_s1_writedata),          //                                                        .writedata
		.key_s1_chipselect                                             (mm_interconnect_1_key_s1_chipselect),         //                                                        .chipselect
		.ledr_s1_address                                               (mm_interconnect_1_ledr_s1_address),           //                                                 ledr_s1.address
		.ledr_s1_write                                                 (mm_interconnect_1_ledr_s1_write),             //                                                        .write
		.ledr_s1_readdata                                              (mm_interconnect_1_ledr_s1_readdata),          //                                                        .readdata
		.ledr_s1_writedata                                             (mm_interconnect_1_ledr_s1_writedata),         //                                                        .writedata
		.ledr_s1_chipselect                                            (mm_interconnect_1_ledr_s1_chipselect),        //                                                        .chipselect
		.sd_clk_s1_address                                             (mm_interconnect_1_sd_clk_s1_address),         //                                               sd_clk_s1.address
		.sd_clk_s1_write                                               (mm_interconnect_1_sd_clk_s1_write),           //                                                        .write
		.sd_clk_s1_readdata                                            (mm_interconnect_1_sd_clk_s1_readdata),        //                                                        .readdata
		.sd_clk_s1_writedata                                           (mm_interconnect_1_sd_clk_s1_writedata),       //                                                        .writedata
		.sd_clk_s1_chipselect                                          (mm_interconnect_1_sd_clk_s1_chipselect),      //                                                        .chipselect
		.sd_cmd_s1_address                                             (mm_interconnect_1_sd_cmd_s1_address),         //                                               sd_cmd_s1.address
		.sd_cmd_s1_write                                               (mm_interconnect_1_sd_cmd_s1_write),           //                                                        .write
		.sd_cmd_s1_readdata                                            (mm_interconnect_1_sd_cmd_s1_readdata),        //                                                        .readdata
		.sd_cmd_s1_writedata                                           (mm_interconnect_1_sd_cmd_s1_writedata),       //                                                        .writedata
		.sd_cmd_s1_chipselect                                          (mm_interconnect_1_sd_cmd_s1_chipselect),      //                                                        .chipselect
		.sd_dat_s1_address                                             (mm_interconnect_1_sd_dat_s1_address),         //                                               sd_dat_s1.address
		.sd_dat_s1_write                                               (mm_interconnect_1_sd_dat_s1_write),           //                                                        .write
		.sd_dat_s1_readdata                                            (mm_interconnect_1_sd_dat_s1_readdata),        //                                                        .readdata
		.sd_dat_s1_writedata                                           (mm_interconnect_1_sd_dat_s1_writedata),       //                                                        .writedata
		.sd_dat_s1_chipselect                                          (mm_interconnect_1_sd_dat_s1_chipselect),      //                                                        .chipselect
		.timer_1_s1_address                                            (mm_interconnect_1_timer_1_s1_address),        //                                              timer_1_s1.address
		.timer_1_s1_write                                              (mm_interconnect_1_timer_1_s1_write),          //                                                        .write
		.timer_1_s1_readdata                                           (mm_interconnect_1_timer_1_s1_readdata),       //                                                        .readdata
		.timer_1_s1_writedata                                          (mm_interconnect_1_timer_1_s1_writedata),      //                                                        .writedata
		.timer_1_s1_chipselect                                         (mm_interconnect_1_timer_1_s1_chipselect)      //                                                        .chipselect
	);

	DE0_CV_system_irq_mapper irq_mapper (
		.clk           (pll_100_outclk0_clk),            //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (cpu_d_irq_irq)                   //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (pll_100_outclk0_clk),                //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (pll_100_outclk0_clk),                //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (pll_100_outclk0_clk),                //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_003 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (pll_100_outclk0_clk),                //         sender_clk.clk
		.receiver_reset (rst_controller_003_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_003_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (pll_100_outclk0_clk),                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_100_outclk0_clk),                //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
